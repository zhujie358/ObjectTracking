////////////////////////////////////////////////////////////////////////////////////////////
// File:   kalman.v
// Author: B. Brown, T. Dotsikas
// About:  Hardware implementation of Kalman filter update equations.
////////////////////////////////////////////////////////////////////////////////////////////

module kalman #(
	parameter COLOR_WIDTH = 10,
	parameter DISP_WIDTH  = 11
)(


);


endmodule